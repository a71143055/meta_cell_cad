module meta_top();
  // cell (0, 0)
  wire cell_0_0_out;
  // cell (1, 0)
  wire cell_1_0_out;
  // cell (2, 0)
  wire cell_2_0_out;
  // cell (3, 0)
  wire cell_3_0_out;
  // cell (4, 0)
  wire cell_4_0_out;
  // cell (5, 0)
  wire cell_5_0_out;
  // cell (6, 0)
  wire cell_6_0_out;
  // cell (7, 0)
  wire cell_7_0_out;
  // cell (8, 0)
  wire cell_8_0_out;
  // cell (9, 0)
  wire cell_9_0_out;
  // cell (10, 0)
  wire cell_10_0_out;
  // cell (11, 0)
  wire cell_11_0_out;
  // cell (0, 1)
  wire cell_0_1_out;
  // cell (1, 1)
  wire cell_1_1_out;
  // cell (2, 1)
  wire cell_2_1_out;
  // cell (3, 1)
  wire cell_3_1_out;
  // cell (4, 1)
  wire cell_4_1_out;
  // cell (5, 1)
  wire cell_5_1_out;
  // cell (6, 1)
  wire cell_6_1_out;
  // cell (7, 1)
  wire cell_7_1_out;
  // cell (8, 1)
  wire cell_8_1_out;
  // cell (9, 1)
  wire cell_9_1_out;
  // cell (10, 1)
  wire cell_10_1_out;
  // cell (11, 1)
  wire cell_11_1_out;
  // cell (0, 2)
  wire cell_0_2_out;
  // cell (1, 2)
  wire cell_1_2_out;
  // cell (2, 2)
  wire cell_2_2_out;
  // cell (3, 2)
  wire cell_3_2_out;
  // cell (4, 2)
  wire cell_4_2_out;
  // cell (5, 2)
  wire cell_5_2_out;
  // cell (6, 2)
  wire cell_6_2_out;
  // cell (7, 2)
  wire cell_7_2_out;
  // cell (8, 2)
  wire cell_8_2_out;
  // cell (9, 2)
  wire cell_9_2_out;
  // cell (10, 2)
  wire cell_10_2_out;
  // cell (11, 2)
  wire cell_11_2_out;
  // cell (0, 3)
  wire cell_0_3_out;
  // cell (1, 3)
  wire cell_1_3_out;
  // cell (2, 3)
  wire cell_2_3_out;
  // cell (3, 3)
  wire cell_3_3_out;
  // cell (4, 3)
  wire cell_4_3_out;
  // cell (5, 3)
  wire cell_5_3_out;
  // cell (6, 3)
  wire cell_6_3_out;
  // cell (7, 3)
  wire cell_7_3_out;
  // cell (8, 3)
  wire cell_8_3_out;
  // cell (9, 3)
  wire cell_9_3_out;
  // cell (10, 3)
  wire cell_10_3_out;
  // cell (11, 3)
  wire cell_11_3_out;
  // cell (0, 4)
  wire cell_0_4_out;
  // cell (1, 4)
  wire cell_1_4_out;
  // cell (2, 4)
  wire cell_2_4_out;
  // cell (3, 4)
  wire cell_3_4_out;
  // cell (4, 4)
  wire cell_4_4_out;
  // cell (5, 4)
  wire cell_5_4_out;
  // cell (6, 4)
  wire cell_6_4_out;
  // cell (7, 4)
  wire cell_7_4_out;
  // cell (8, 4)
  wire cell_8_4_out;
  // cell (9, 4)
  wire cell_9_4_out;
  // cell (10, 4)
  wire cell_10_4_out;
  // cell (11, 4)
  wire cell_11_4_out;
  // cell (0, 5)
  wire cell_0_5_out;
  // cell (1, 5)
  wire cell_1_5_out;
  // cell (2, 5)
  wire cell_2_5_out;
  // cell (3, 5)
  wire cell_3_5_out;
  // cell (4, 5)
  wire cell_4_5_out;
  // cell (5, 5)
  wire cell_5_5_out;
  // cell (6, 5)
  wire cell_6_5_out;
  // cell (7, 5)
  wire cell_7_5_out;
  // cell (8, 5)
  wire cell_8_5_out;
  // cell (9, 5)
  wire cell_9_5_out;
  // cell (10, 5)
  wire cell_10_5_out;
  // cell (11, 5)
  wire cell_11_5_out;
  // cell (0, 6)
  wire cell_0_6_out;
  // cell (1, 6)
  wire cell_1_6_out;
  // cell (2, 6)
  wire cell_2_6_out;
  // cell (3, 6)
  wire cell_3_6_out;
  // cell (4, 6)
  wire cell_4_6_out;
  // cell (5, 6)
  wire cell_5_6_out;
  // cell (6, 6)
  wire cell_6_6_out;
  // cell (7, 6)
  wire cell_7_6_out;
  // cell (8, 6)
  wire cell_8_6_out;
  // cell (9, 6)
  wire cell_9_6_out;
  // cell (10, 6)
  wire cell_10_6_out;
  // cell (11, 6)
  wire cell_11_6_out;
  // cell (0, 7)
  wire cell_0_7_out;
  // cell (1, 7)
  wire cell_1_7_out;
  // cell (2, 7)
  wire cell_2_7_out;
  // cell (3, 7)
  wire cell_3_7_out;
  // cell (4, 7)
  wire cell_4_7_out;
  // cell (5, 7)
  wire cell_5_7_out;
  // cell (6, 7)
  wire cell_6_7_out;
  // cell (7, 7)
  wire cell_7_7_out;
  // cell (8, 7)
  wire cell_8_7_out;
  // cell (9, 7)
  wire cell_9_7_out;
  // cell (10, 7)
  wire cell_10_7_out;
  // cell (11, 7)
  wire cell_11_7_out;
  // cell (0, 8)
  wire cell_0_8_out;
  // cell (1, 8)
  wire cell_1_8_out;
  // cell (2, 8)
  wire cell_2_8_out;
  // cell (3, 8)
  wire cell_3_8_out;
  // cell (4, 8)
  wire cell_4_8_out;
  // cell (5, 8)
  wire cell_5_8_out;
  // cell (6, 8)
  wire cell_6_8_out;
  // cell (7, 8)
  wire cell_7_8_out;
  // cell (8, 8)
  wire cell_8_8_out;
  // cell (9, 8)
  wire cell_9_8_out;
  // cell (10, 8)
  wire cell_10_8_out;
  // cell (11, 8)
  wire cell_11_8_out;
  // cell (0, 9)
  wire cell_0_9_out;
  // cell (1, 9)
  wire cell_1_9_out;
  // cell (2, 9)
  wire cell_2_9_out;
  // cell (3, 9)
  wire cell_3_9_out;
  // cell (4, 9)
  wire cell_4_9_out;
  // cell (5, 9)
  wire cell_5_9_out;
  // cell (6, 9)
  wire cell_6_9_out;
  // cell (7, 9)
  wire cell_7_9_out;
  // cell (8, 9)
  wire cell_8_9_out;
  // cell (9, 9)
  wire cell_9_9_out;
  // cell (10, 9)
  wire cell_10_9_out;
  // cell (11, 9)
  wire cell_11_9_out;
  // cell (0, 10)
  wire cell_0_10_out;
  // cell (1, 10)
  wire cell_1_10_out;
  // cell (2, 10)
  wire cell_2_10_out;
  // cell (3, 10)
  wire cell_3_10_out;
  // cell (4, 10)
  wire cell_4_10_out;
  // cell (5, 10)
  wire cell_5_10_out;
  // cell (6, 10)
  wire cell_6_10_out;
  // cell (7, 10)
  wire cell_7_10_out;
  // cell (8, 10)
  wire cell_8_10_out;
  // cell (9, 10)
  wire cell_9_10_out;
  // cell (10, 10)
  wire cell_10_10_out;
  // cell (11, 10)
  wire cell_11_10_out;
  // cell (0, 11)
  wire cell_0_11_out;
  // cell (1, 11)
  wire cell_1_11_out;
  // cell (2, 11)
  wire cell_2_11_out;
  // cell (3, 11)
  wire cell_3_11_out;
  // cell (4, 11)
  wire cell_4_11_out;
  // cell (5, 11)
  wire cell_5_11_out;
  // cell (6, 11)
  wire cell_6_11_out;
  // cell (7, 11)
  wire cell_7_11_out;
  // cell (8, 11)
  wire cell_8_11_out;
  // cell (9, 11)
  wire cell_9_11_out;
  // cell (10, 11)
  wire cell_10_11_out;
  // cell (11, 11)
  wire cell_11_11_out;
  // (0, 0) -> (1, 0) (out)
  assign cell_1_0_out = cell_0_0_out;
  // (0, 0) -> (0, 1) (out)
  assign cell_0_1_out = cell_0_0_out;
  // (1, 0) -> (2, 0) (out)
  assign cell_2_0_out = cell_1_0_out;
  // (1, 0) -> (0, 0) (out)
  assign cell_0_0_out = cell_1_0_out;
  // (1, 0) -> (1, 1) (out)
  assign cell_1_1_out = cell_1_0_out;
  // (2, 0) -> (3, 0) (out)
  assign cell_3_0_out = cell_2_0_out;
  // (2, 0) -> (1, 0) (out)
  assign cell_1_0_out = cell_2_0_out;
  // (2, 0) -> (2, 1) (out)
  assign cell_2_1_out = cell_2_0_out;
  // (3, 0) -> (4, 0) (out)
  assign cell_4_0_out = cell_3_0_out;
  // (3, 0) -> (2, 0) (out)
  assign cell_2_0_out = cell_3_0_out;
  // (3, 0) -> (3, 1) (out)
  assign cell_3_1_out = cell_3_0_out;
  // (4, 0) -> (5, 0) (out)
  assign cell_5_0_out = cell_4_0_out;
  // (4, 0) -> (3, 0) (out)
  assign cell_3_0_out = cell_4_0_out;
  // (4, 0) -> (4, 1) (out)
  assign cell_4_1_out = cell_4_0_out;
  // (5, 0) -> (6, 0) (out)
  assign cell_6_0_out = cell_5_0_out;
  // (5, 0) -> (4, 0) (out)
  assign cell_4_0_out = cell_5_0_out;
  // (5, 0) -> (5, 1) (out)
  assign cell_5_1_out = cell_5_0_out;
  // (6, 0) -> (7, 0) (out)
  assign cell_7_0_out = cell_6_0_out;
  // (6, 0) -> (5, 0) (out)
  assign cell_5_0_out = cell_6_0_out;
  // (6, 0) -> (6, 1) (out)
  assign cell_6_1_out = cell_6_0_out;
  // (7, 0) -> (8, 0) (out)
  assign cell_8_0_out = cell_7_0_out;
  // (7, 0) -> (6, 0) (out)
  assign cell_6_0_out = cell_7_0_out;
  // (7, 0) -> (7, 1) (out)
  assign cell_7_1_out = cell_7_0_out;
  // (8, 0) -> (9, 0) (out)
  assign cell_9_0_out = cell_8_0_out;
  // (8, 0) -> (7, 0) (out)
  assign cell_7_0_out = cell_8_0_out;
  // (8, 0) -> (8, 1) (out)
  assign cell_8_1_out = cell_8_0_out;
  // (9, 0) -> (10, 0) (out)
  assign cell_10_0_out = cell_9_0_out;
  // (9, 0) -> (8, 0) (out)
  assign cell_8_0_out = cell_9_0_out;
  // (9, 0) -> (9, 1) (out)
  assign cell_9_1_out = cell_9_0_out;
  // (10, 0) -> (11, 0) (out)
  assign cell_11_0_out = cell_10_0_out;
  // (10, 0) -> (9, 0) (out)
  assign cell_9_0_out = cell_10_0_out;
  // (10, 0) -> (10, 1) (out)
  assign cell_10_1_out = cell_10_0_out;
  // (11, 0) -> (10, 0) (out)
  assign cell_10_0_out = cell_11_0_out;
  // (11, 0) -> (11, 1) (out)
  assign cell_11_1_out = cell_11_0_out;
  // (0, 1) -> (1, 1) (out)
  assign cell_1_1_out = cell_0_1_out;
  // (0, 1) -> (0, 2) (out)
  assign cell_0_2_out = cell_0_1_out;
  // (0, 1) -> (0, 0) (out)
  assign cell_0_0_out = cell_0_1_out;
  // (1, 1) -> (2, 1) (out)
  assign cell_2_1_out = cell_1_1_out;
  // (1, 1) -> (0, 1) (out)
  assign cell_0_1_out = cell_1_1_out;
  // (1, 1) -> (1, 2) (out)
  assign cell_1_2_out = cell_1_1_out;
  // (1, 1) -> (1, 0) (out)
  assign cell_1_0_out = cell_1_1_out;
  // (2, 1) -> (3, 1) (out)
  assign cell_3_1_out = cell_2_1_out;
  // (2, 1) -> (1, 1) (out)
  assign cell_1_1_out = cell_2_1_out;
  // (2, 1) -> (2, 2) (out)
  assign cell_2_2_out = cell_2_1_out;
  // (2, 1) -> (2, 0) (out)
  assign cell_2_0_out = cell_2_1_out;
  // (3, 1) -> (4, 1) (out)
  assign cell_4_1_out = cell_3_1_out;
  // (3, 1) -> (2, 1) (out)
  assign cell_2_1_out = cell_3_1_out;
  // (3, 1) -> (3, 2) (out)
  assign cell_3_2_out = cell_3_1_out;
  // (3, 1) -> (3, 0) (out)
  assign cell_3_0_out = cell_3_1_out;
  // (4, 1) -> (5, 1) (out)
  assign cell_5_1_out = cell_4_1_out;
  // (4, 1) -> (3, 1) (out)
  assign cell_3_1_out = cell_4_1_out;
  // (4, 1) -> (4, 2) (out)
  assign cell_4_2_out = cell_4_1_out;
  // (4, 1) -> (4, 0) (out)
  assign cell_4_0_out = cell_4_1_out;
  // (5, 1) -> (6, 1) (out)
  assign cell_6_1_out = cell_5_1_out;
  // (5, 1) -> (4, 1) (out)
  assign cell_4_1_out = cell_5_1_out;
  // (5, 1) -> (5, 2) (out)
  assign cell_5_2_out = cell_5_1_out;
  // (5, 1) -> (5, 0) (out)
  assign cell_5_0_out = cell_5_1_out;
  // (6, 1) -> (7, 1) (out)
  assign cell_7_1_out = cell_6_1_out;
  // (6, 1) -> (5, 1) (out)
  assign cell_5_1_out = cell_6_1_out;
  // (6, 1) -> (6, 2) (out)
  assign cell_6_2_out = cell_6_1_out;
  // (6, 1) -> (6, 0) (out)
  assign cell_6_0_out = cell_6_1_out;
  // (7, 1) -> (8, 1) (out)
  assign cell_8_1_out = cell_7_1_out;
  // (7, 1) -> (6, 1) (out)
  assign cell_6_1_out = cell_7_1_out;
  // (7, 1) -> (7, 2) (out)
  assign cell_7_2_out = cell_7_1_out;
  // (7, 1) -> (7, 0) (out)
  assign cell_7_0_out = cell_7_1_out;
  // (8, 1) -> (9, 1) (out)
  assign cell_9_1_out = cell_8_1_out;
  // (8, 1) -> (7, 1) (out)
  assign cell_7_1_out = cell_8_1_out;
  // (8, 1) -> (8, 2) (out)
  assign cell_8_2_out = cell_8_1_out;
  // (8, 1) -> (8, 0) (out)
  assign cell_8_0_out = cell_8_1_out;
  // (9, 1) -> (10, 1) (out)
  assign cell_10_1_out = cell_9_1_out;
  // (9, 1) -> (8, 1) (out)
  assign cell_8_1_out = cell_9_1_out;
  // (9, 1) -> (9, 2) (out)
  assign cell_9_2_out = cell_9_1_out;
  // (9, 1) -> (9, 0) (out)
  assign cell_9_0_out = cell_9_1_out;
  // (10, 1) -> (11, 1) (out)
  assign cell_11_1_out = cell_10_1_out;
  // (10, 1) -> (9, 1) (out)
  assign cell_9_1_out = cell_10_1_out;
  // (10, 1) -> (10, 2) (out)
  assign cell_10_2_out = cell_10_1_out;
  // (10, 1) -> (10, 0) (out)
  assign cell_10_0_out = cell_10_1_out;
  // (11, 1) -> (10, 1) (out)
  assign cell_10_1_out = cell_11_1_out;
  // (11, 1) -> (11, 2) (out)
  assign cell_11_2_out = cell_11_1_out;
  // (11, 1) -> (11, 0) (out)
  assign cell_11_0_out = cell_11_1_out;
  // (0, 2) -> (1, 2) (out)
  assign cell_1_2_out = cell_0_2_out;
  // (0, 2) -> (0, 3) (out)
  assign cell_0_3_out = cell_0_2_out;
  // (0, 2) -> (0, 1) (out)
  assign cell_0_1_out = cell_0_2_out;
  // (1, 2) -> (2, 2) (out)
  assign cell_2_2_out = cell_1_2_out;
  // (1, 2) -> (0, 2) (out)
  assign cell_0_2_out = cell_1_2_out;
  // (1, 2) -> (1, 3) (out)
  assign cell_1_3_out = cell_1_2_out;
  // (1, 2) -> (1, 1) (out)
  assign cell_1_1_out = cell_1_2_out;
  // (2, 2) -> (3, 2) (out)
  assign cell_3_2_out = cell_2_2_out;
  // (2, 2) -> (1, 2) (out)
  assign cell_1_2_out = cell_2_2_out;
  // (2, 2) -> (2, 3) (out)
  assign cell_2_3_out = cell_2_2_out;
  // (2, 2) -> (2, 1) (out)
  assign cell_2_1_out = cell_2_2_out;
  // (3, 2) -> (4, 2) (out)
  assign cell_4_2_out = cell_3_2_out;
  // (3, 2) -> (2, 2) (out)
  assign cell_2_2_out = cell_3_2_out;
  // (3, 2) -> (3, 3) (out)
  assign cell_3_3_out = cell_3_2_out;
  // (3, 2) -> (3, 1) (out)
  assign cell_3_1_out = cell_3_2_out;
  // (4, 2) -> (5, 2) (out)
  assign cell_5_2_out = cell_4_2_out;
  // (4, 2) -> (3, 2) (out)
  assign cell_3_2_out = cell_4_2_out;
  // (4, 2) -> (4, 3) (out)
  assign cell_4_3_out = cell_4_2_out;
  // (4, 2) -> (4, 1) (out)
  assign cell_4_1_out = cell_4_2_out;
  // (5, 2) -> (6, 2) (out)
  assign cell_6_2_out = cell_5_2_out;
  // (5, 2) -> (4, 2) (out)
  assign cell_4_2_out = cell_5_2_out;
  // (5, 2) -> (5, 3) (out)
  assign cell_5_3_out = cell_5_2_out;
  // (5, 2) -> (5, 1) (out)
  assign cell_5_1_out = cell_5_2_out;
  // (6, 2) -> (7, 2) (out)
  assign cell_7_2_out = cell_6_2_out;
  // (6, 2) -> (5, 2) (out)
  assign cell_5_2_out = cell_6_2_out;
  // (6, 2) -> (6, 3) (out)
  assign cell_6_3_out = cell_6_2_out;
  // (6, 2) -> (6, 1) (out)
  assign cell_6_1_out = cell_6_2_out;
  // (7, 2) -> (8, 2) (out)
  assign cell_8_2_out = cell_7_2_out;
  // (7, 2) -> (6, 2) (out)
  assign cell_6_2_out = cell_7_2_out;
  // (7, 2) -> (7, 3) (out)
  assign cell_7_3_out = cell_7_2_out;
  // (7, 2) -> (7, 1) (out)
  assign cell_7_1_out = cell_7_2_out;
  // (8, 2) -> (9, 2) (out)
  assign cell_9_2_out = cell_8_2_out;
  // (8, 2) -> (7, 2) (out)
  assign cell_7_2_out = cell_8_2_out;
  // (8, 2) -> (8, 3) (out)
  assign cell_8_3_out = cell_8_2_out;
  // (8, 2) -> (8, 1) (out)
  assign cell_8_1_out = cell_8_2_out;
  // (9, 2) -> (10, 2) (out)
  assign cell_10_2_out = cell_9_2_out;
  // (9, 2) -> (8, 2) (out)
  assign cell_8_2_out = cell_9_2_out;
  // (9, 2) -> (9, 3) (out)
  assign cell_9_3_out = cell_9_2_out;
  // (9, 2) -> (9, 1) (out)
  assign cell_9_1_out = cell_9_2_out;
  // (10, 2) -> (11, 2) (out)
  assign cell_11_2_out = cell_10_2_out;
  // (10, 2) -> (9, 2) (out)
  assign cell_9_2_out = cell_10_2_out;
  // (10, 2) -> (10, 3) (out)
  assign cell_10_3_out = cell_10_2_out;
  // (10, 2) -> (10, 1) (out)
  assign cell_10_1_out = cell_10_2_out;
  // (11, 2) -> (10, 2) (out)
  assign cell_10_2_out = cell_11_2_out;
  // (11, 2) -> (11, 3) (out)
  assign cell_11_3_out = cell_11_2_out;
  // (11, 2) -> (11, 1) (out)
  assign cell_11_1_out = cell_11_2_out;
  // (0, 3) -> (1, 3) (out)
  assign cell_1_3_out = cell_0_3_out;
  // (0, 3) -> (0, 4) (out)
  assign cell_0_4_out = cell_0_3_out;
  // (0, 3) -> (0, 2) (out)
  assign cell_0_2_out = cell_0_3_out;
  // (1, 3) -> (2, 3) (out)
  assign cell_2_3_out = cell_1_3_out;
  // (1, 3) -> (0, 3) (out)
  assign cell_0_3_out = cell_1_3_out;
  // (1, 3) -> (1, 4) (out)
  assign cell_1_4_out = cell_1_3_out;
  // (1, 3) -> (1, 2) (out)
  assign cell_1_2_out = cell_1_3_out;
  // (2, 3) -> (3, 3) (out)
  assign cell_3_3_out = cell_2_3_out;
  // (2, 3) -> (1, 3) (out)
  assign cell_1_3_out = cell_2_3_out;
  // (2, 3) -> (2, 4) (out)
  assign cell_2_4_out = cell_2_3_out;
  // (2, 3) -> (2, 2) (out)
  assign cell_2_2_out = cell_2_3_out;
  // (3, 3) -> (4, 3) (out)
  assign cell_4_3_out = cell_3_3_out;
  // (3, 3) -> (2, 3) (out)
  assign cell_2_3_out = cell_3_3_out;
  // (3, 3) -> (3, 4) (out)
  assign cell_3_4_out = cell_3_3_out;
  // (3, 3) -> (3, 2) (out)
  assign cell_3_2_out = cell_3_3_out;
  // (4, 3) -> (5, 3) (out)
  assign cell_5_3_out = cell_4_3_out;
  // (4, 3) -> (3, 3) (out)
  assign cell_3_3_out = cell_4_3_out;
  // (4, 3) -> (4, 4) (out)
  assign cell_4_4_out = cell_4_3_out;
  // (4, 3) -> (4, 2) (out)
  assign cell_4_2_out = cell_4_3_out;
  // (5, 3) -> (6, 3) (out)
  assign cell_6_3_out = cell_5_3_out;
  // (5, 3) -> (4, 3) (out)
  assign cell_4_3_out = cell_5_3_out;
  // (5, 3) -> (5, 4) (out)
  assign cell_5_4_out = cell_5_3_out;
  // (5, 3) -> (5, 2) (out)
  assign cell_5_2_out = cell_5_3_out;
  // (6, 3) -> (7, 3) (out)
  assign cell_7_3_out = cell_6_3_out;
  // (6, 3) -> (5, 3) (out)
  assign cell_5_3_out = cell_6_3_out;
  // (6, 3) -> (6, 4) (out)
  assign cell_6_4_out = cell_6_3_out;
  // (6, 3) -> (6, 2) (out)
  assign cell_6_2_out = cell_6_3_out;
  // (7, 3) -> (8, 3) (out)
  assign cell_8_3_out = cell_7_3_out;
  // (7, 3) -> (6, 3) (out)
  assign cell_6_3_out = cell_7_3_out;
  // (7, 3) -> (7, 4) (out)
  assign cell_7_4_out = cell_7_3_out;
  // (7, 3) -> (7, 2) (out)
  assign cell_7_2_out = cell_7_3_out;
  // (8, 3) -> (9, 3) (out)
  assign cell_9_3_out = cell_8_3_out;
  // (8, 3) -> (7, 3) (out)
  assign cell_7_3_out = cell_8_3_out;
  // (8, 3) -> (8, 4) (out)
  assign cell_8_4_out = cell_8_3_out;
  // (8, 3) -> (8, 2) (out)
  assign cell_8_2_out = cell_8_3_out;
  // (9, 3) -> (10, 3) (out)
  assign cell_10_3_out = cell_9_3_out;
  // (9, 3) -> (8, 3) (out)
  assign cell_8_3_out = cell_9_3_out;
  // (9, 3) -> (9, 4) (out)
  assign cell_9_4_out = cell_9_3_out;
  // (9, 3) -> (9, 2) (out)
  assign cell_9_2_out = cell_9_3_out;
  // (10, 3) -> (11, 3) (out)
  assign cell_11_3_out = cell_10_3_out;
  // (10, 3) -> (9, 3) (out)
  assign cell_9_3_out = cell_10_3_out;
  // (10, 3) -> (10, 4) (out)
  assign cell_10_4_out = cell_10_3_out;
  // (10, 3) -> (10, 2) (out)
  assign cell_10_2_out = cell_10_3_out;
  // (11, 3) -> (10, 3) (out)
  assign cell_10_3_out = cell_11_3_out;
  // (11, 3) -> (11, 4) (out)
  assign cell_11_4_out = cell_11_3_out;
  // (11, 3) -> (11, 2) (out)
  assign cell_11_2_out = cell_11_3_out;
  // (0, 4) -> (1, 4) (out)
  assign cell_1_4_out = cell_0_4_out;
  // (0, 4) -> (0, 5) (out)
  assign cell_0_5_out = cell_0_4_out;
  // (0, 4) -> (0, 3) (out)
  assign cell_0_3_out = cell_0_4_out;
  // (1, 4) -> (2, 4) (out)
  assign cell_2_4_out = cell_1_4_out;
  // (1, 4) -> (0, 4) (out)
  assign cell_0_4_out = cell_1_4_out;
  // (1, 4) -> (1, 5) (out)
  assign cell_1_5_out = cell_1_4_out;
  // (1, 4) -> (1, 3) (out)
  assign cell_1_3_out = cell_1_4_out;
  // (2, 4) -> (3, 4) (out)
  assign cell_3_4_out = cell_2_4_out;
  // (2, 4) -> (1, 4) (out)
  assign cell_1_4_out = cell_2_4_out;
  // (2, 4) -> (2, 5) (out)
  assign cell_2_5_out = cell_2_4_out;
  // (2, 4) -> (2, 3) (out)
  assign cell_2_3_out = cell_2_4_out;
  // (3, 4) -> (4, 4) (out)
  assign cell_4_4_out = cell_3_4_out;
  // (3, 4) -> (2, 4) (out)
  assign cell_2_4_out = cell_3_4_out;
  // (3, 4) -> (3, 5) (out)
  assign cell_3_5_out = cell_3_4_out;
  // (3, 4) -> (3, 3) (out)
  assign cell_3_3_out = cell_3_4_out;
  // (4, 4) -> (5, 4) (out)
  assign cell_5_4_out = cell_4_4_out;
  // (4, 4) -> (3, 4) (out)
  assign cell_3_4_out = cell_4_4_out;
  // (4, 4) -> (4, 5) (out)
  assign cell_4_5_out = cell_4_4_out;
  // (4, 4) -> (4, 3) (out)
  assign cell_4_3_out = cell_4_4_out;
  // (5, 4) -> (6, 4) (out)
  assign cell_6_4_out = cell_5_4_out;
  // (5, 4) -> (4, 4) (out)
  assign cell_4_4_out = cell_5_4_out;
  // (5, 4) -> (5, 5) (out)
  assign cell_5_5_out = cell_5_4_out;
  // (5, 4) -> (5, 3) (out)
  assign cell_5_3_out = cell_5_4_out;
  // (6, 4) -> (7, 4) (out)
  assign cell_7_4_out = cell_6_4_out;
  // (6, 4) -> (5, 4) (out)
  assign cell_5_4_out = cell_6_4_out;
  // (6, 4) -> (6, 5) (out)
  assign cell_6_5_out = cell_6_4_out;
  // (6, 4) -> (6, 3) (out)
  assign cell_6_3_out = cell_6_4_out;
  // (7, 4) -> (8, 4) (out)
  assign cell_8_4_out = cell_7_4_out;
  // (7, 4) -> (6, 4) (out)
  assign cell_6_4_out = cell_7_4_out;
  // (7, 4) -> (7, 5) (out)
  assign cell_7_5_out = cell_7_4_out;
  // (7, 4) -> (7, 3) (out)
  assign cell_7_3_out = cell_7_4_out;
  // (8, 4) -> (9, 4) (out)
  assign cell_9_4_out = cell_8_4_out;
  // (8, 4) -> (7, 4) (out)
  assign cell_7_4_out = cell_8_4_out;
  // (8, 4) -> (8, 5) (out)
  assign cell_8_5_out = cell_8_4_out;
  // (8, 4) -> (8, 3) (out)
  assign cell_8_3_out = cell_8_4_out;
  // (9, 4) -> (10, 4) (out)
  assign cell_10_4_out = cell_9_4_out;
  // (9, 4) -> (8, 4) (out)
  assign cell_8_4_out = cell_9_4_out;
  // (9, 4) -> (9, 5) (out)
  assign cell_9_5_out = cell_9_4_out;
  // (9, 4) -> (9, 3) (out)
  assign cell_9_3_out = cell_9_4_out;
  // (10, 4) -> (11, 4) (out)
  assign cell_11_4_out = cell_10_4_out;
  // (10, 4) -> (9, 4) (out)
  assign cell_9_4_out = cell_10_4_out;
  // (10, 4) -> (10, 5) (out)
  assign cell_10_5_out = cell_10_4_out;
  // (10, 4) -> (10, 3) (out)
  assign cell_10_3_out = cell_10_4_out;
  // (11, 4) -> (10, 4) (out)
  assign cell_10_4_out = cell_11_4_out;
  // (11, 4) -> (11, 5) (out)
  assign cell_11_5_out = cell_11_4_out;
  // (11, 4) -> (11, 3) (out)
  assign cell_11_3_out = cell_11_4_out;
  // (0, 5) -> (1, 5) (out)
  assign cell_1_5_out = cell_0_5_out;
  // (0, 5) -> (0, 6) (out)
  assign cell_0_6_out = cell_0_5_out;
  // (0, 5) -> (0, 4) (out)
  assign cell_0_4_out = cell_0_5_out;
  // (1, 5) -> (2, 5) (out)
  assign cell_2_5_out = cell_1_5_out;
  // (1, 5) -> (0, 5) (out)
  assign cell_0_5_out = cell_1_5_out;
  // (1, 5) -> (1, 6) (out)
  assign cell_1_6_out = cell_1_5_out;
  // (1, 5) -> (1, 4) (out)
  assign cell_1_4_out = cell_1_5_out;
  // (2, 5) -> (3, 5) (out)
  assign cell_3_5_out = cell_2_5_out;
  // (2, 5) -> (1, 5) (out)
  assign cell_1_5_out = cell_2_5_out;
  // (2, 5) -> (2, 6) (out)
  assign cell_2_6_out = cell_2_5_out;
  // (2, 5) -> (2, 4) (out)
  assign cell_2_4_out = cell_2_5_out;
  // (3, 5) -> (4, 5) (out)
  assign cell_4_5_out = cell_3_5_out;
  // (3, 5) -> (2, 5) (out)
  assign cell_2_5_out = cell_3_5_out;
  // (3, 5) -> (3, 6) (out)
  assign cell_3_6_out = cell_3_5_out;
  // (3, 5) -> (3, 4) (out)
  assign cell_3_4_out = cell_3_5_out;
  // (4, 5) -> (5, 5) (out)
  assign cell_5_5_out = cell_4_5_out;
  // (4, 5) -> (3, 5) (out)
  assign cell_3_5_out = cell_4_5_out;
  // (4, 5) -> (4, 6) (out)
  assign cell_4_6_out = cell_4_5_out;
  // (4, 5) -> (4, 4) (out)
  assign cell_4_4_out = cell_4_5_out;
  // (5, 5) -> (6, 5) (out)
  assign cell_6_5_out = cell_5_5_out;
  // (5, 5) -> (4, 5) (out)
  assign cell_4_5_out = cell_5_5_out;
  // (5, 5) -> (5, 6) (out)
  assign cell_5_6_out = cell_5_5_out;
  // (5, 5) -> (5, 4) (out)
  assign cell_5_4_out = cell_5_5_out;
  // (6, 5) -> (7, 5) (out)
  assign cell_7_5_out = cell_6_5_out;
  // (6, 5) -> (5, 5) (out)
  assign cell_5_5_out = cell_6_5_out;
  // (6, 5) -> (6, 6) (out)
  assign cell_6_6_out = cell_6_5_out;
  // (6, 5) -> (6, 4) (out)
  assign cell_6_4_out = cell_6_5_out;
  // (7, 5) -> (8, 5) (out)
  assign cell_8_5_out = cell_7_5_out;
  // (7, 5) -> (6, 5) (out)
  assign cell_6_5_out = cell_7_5_out;
  // (7, 5) -> (7, 6) (out)
  assign cell_7_6_out = cell_7_5_out;
  // (7, 5) -> (7, 4) (out)
  assign cell_7_4_out = cell_7_5_out;
  // (8, 5) -> (9, 5) (out)
  assign cell_9_5_out = cell_8_5_out;
  // (8, 5) -> (7, 5) (out)
  assign cell_7_5_out = cell_8_5_out;
  // (8, 5) -> (8, 6) (out)
  assign cell_8_6_out = cell_8_5_out;
  // (8, 5) -> (8, 4) (out)
  assign cell_8_4_out = cell_8_5_out;
  // (9, 5) -> (10, 5) (out)
  assign cell_10_5_out = cell_9_5_out;
  // (9, 5) -> (8, 5) (out)
  assign cell_8_5_out = cell_9_5_out;
  // (9, 5) -> (9, 6) (out)
  assign cell_9_6_out = cell_9_5_out;
  // (9, 5) -> (9, 4) (out)
  assign cell_9_4_out = cell_9_5_out;
  // (10, 5) -> (11, 5) (out)
  assign cell_11_5_out = cell_10_5_out;
  // (10, 5) -> (9, 5) (out)
  assign cell_9_5_out = cell_10_5_out;
  // (10, 5) -> (10, 6) (out)
  assign cell_10_6_out = cell_10_5_out;
  // (10, 5) -> (10, 4) (out)
  assign cell_10_4_out = cell_10_5_out;
  // (11, 5) -> (10, 5) (out)
  assign cell_10_5_out = cell_11_5_out;
  // (11, 5) -> (11, 6) (out)
  assign cell_11_6_out = cell_11_5_out;
  // (11, 5) -> (11, 4) (out)
  assign cell_11_4_out = cell_11_5_out;
  // (0, 6) -> (1, 6) (out)
  assign cell_1_6_out = cell_0_6_out;
  // (0, 6) -> (0, 7) (out)
  assign cell_0_7_out = cell_0_6_out;
  // (0, 6) -> (0, 5) (out)
  assign cell_0_5_out = cell_0_6_out;
  // (1, 6) -> (2, 6) (out)
  assign cell_2_6_out = cell_1_6_out;
  // (1, 6) -> (0, 6) (out)
  assign cell_0_6_out = cell_1_6_out;
  // (1, 6) -> (1, 7) (out)
  assign cell_1_7_out = cell_1_6_out;
  // (1, 6) -> (1, 5) (out)
  assign cell_1_5_out = cell_1_6_out;
  // (2, 6) -> (3, 6) (out)
  assign cell_3_6_out = cell_2_6_out;
  // (2, 6) -> (1, 6) (out)
  assign cell_1_6_out = cell_2_6_out;
  // (2, 6) -> (2, 7) (out)
  assign cell_2_7_out = cell_2_6_out;
  // (2, 6) -> (2, 5) (out)
  assign cell_2_5_out = cell_2_6_out;
  // (3, 6) -> (4, 6) (out)
  assign cell_4_6_out = cell_3_6_out;
  // (3, 6) -> (2, 6) (out)
  assign cell_2_6_out = cell_3_6_out;
  // (3, 6) -> (3, 7) (out)
  assign cell_3_7_out = cell_3_6_out;
  // (3, 6) -> (3, 5) (out)
  assign cell_3_5_out = cell_3_6_out;
  // (4, 6) -> (5, 6) (out)
  assign cell_5_6_out = cell_4_6_out;
  // (4, 6) -> (3, 6) (out)
  assign cell_3_6_out = cell_4_6_out;
  // (4, 6) -> (4, 7) (out)
  assign cell_4_7_out = cell_4_6_out;
  // (4, 6) -> (4, 5) (out)
  assign cell_4_5_out = cell_4_6_out;
  // (5, 6) -> (6, 6) (out)
  assign cell_6_6_out = cell_5_6_out;
  // (5, 6) -> (4, 6) (out)
  assign cell_4_6_out = cell_5_6_out;
  // (5, 6) -> (5, 7) (out)
  assign cell_5_7_out = cell_5_6_out;
  // (5, 6) -> (5, 5) (out)
  assign cell_5_5_out = cell_5_6_out;
  // (6, 6) -> (7, 6) (out)
  assign cell_7_6_out = cell_6_6_out;
  // (6, 6) -> (5, 6) (out)
  assign cell_5_6_out = cell_6_6_out;
  // (6, 6) -> (6, 7) (out)
  assign cell_6_7_out = cell_6_6_out;
  // (6, 6) -> (6, 5) (out)
  assign cell_6_5_out = cell_6_6_out;
  // (7, 6) -> (8, 6) (out)
  assign cell_8_6_out = cell_7_6_out;
  // (7, 6) -> (6, 6) (out)
  assign cell_6_6_out = cell_7_6_out;
  // (7, 6) -> (7, 7) (out)
  assign cell_7_7_out = cell_7_6_out;
  // (7, 6) -> (7, 5) (out)
  assign cell_7_5_out = cell_7_6_out;
  // (8, 6) -> (9, 6) (out)
  assign cell_9_6_out = cell_8_6_out;
  // (8, 6) -> (7, 6) (out)
  assign cell_7_6_out = cell_8_6_out;
  // (8, 6) -> (8, 7) (out)
  assign cell_8_7_out = cell_8_6_out;
  // (8, 6) -> (8, 5) (out)
  assign cell_8_5_out = cell_8_6_out;
  // (9, 6) -> (10, 6) (out)
  assign cell_10_6_out = cell_9_6_out;
  // (9, 6) -> (8, 6) (out)
  assign cell_8_6_out = cell_9_6_out;
  // (9, 6) -> (9, 7) (out)
  assign cell_9_7_out = cell_9_6_out;
  // (9, 6) -> (9, 5) (out)
  assign cell_9_5_out = cell_9_6_out;
  // (10, 6) -> (11, 6) (out)
  assign cell_11_6_out = cell_10_6_out;
  // (10, 6) -> (9, 6) (out)
  assign cell_9_6_out = cell_10_6_out;
  // (10, 6) -> (10, 7) (out)
  assign cell_10_7_out = cell_10_6_out;
  // (10, 6) -> (10, 5) (out)
  assign cell_10_5_out = cell_10_6_out;
  // (11, 6) -> (10, 6) (out)
  assign cell_10_6_out = cell_11_6_out;
  // (11, 6) -> (11, 7) (out)
  assign cell_11_7_out = cell_11_6_out;
  // (11, 6) -> (11, 5) (out)
  assign cell_11_5_out = cell_11_6_out;
  // (0, 7) -> (1, 7) (out)
  assign cell_1_7_out = cell_0_7_out;
  // (0, 7) -> (0, 8) (out)
  assign cell_0_8_out = cell_0_7_out;
  // (0, 7) -> (0, 6) (out)
  assign cell_0_6_out = cell_0_7_out;
  // (1, 7) -> (2, 7) (out)
  assign cell_2_7_out = cell_1_7_out;
  // (1, 7) -> (0, 7) (out)
  assign cell_0_7_out = cell_1_7_out;
  // (1, 7) -> (1, 8) (out)
  assign cell_1_8_out = cell_1_7_out;
  // (1, 7) -> (1, 6) (out)
  assign cell_1_6_out = cell_1_7_out;
  // (2, 7) -> (3, 7) (out)
  assign cell_3_7_out = cell_2_7_out;
  // (2, 7) -> (1, 7) (out)
  assign cell_1_7_out = cell_2_7_out;
  // (2, 7) -> (2, 8) (out)
  assign cell_2_8_out = cell_2_7_out;
  // (2, 7) -> (2, 6) (out)
  assign cell_2_6_out = cell_2_7_out;
  // (3, 7) -> (4, 7) (out)
  assign cell_4_7_out = cell_3_7_out;
  // (3, 7) -> (2, 7) (out)
  assign cell_2_7_out = cell_3_7_out;
  // (3, 7) -> (3, 8) (out)
  assign cell_3_8_out = cell_3_7_out;
  // (3, 7) -> (3, 6) (out)
  assign cell_3_6_out = cell_3_7_out;
  // (4, 7) -> (5, 7) (out)
  assign cell_5_7_out = cell_4_7_out;
  // (4, 7) -> (3, 7) (out)
  assign cell_3_7_out = cell_4_7_out;
  // (4, 7) -> (4, 8) (out)
  assign cell_4_8_out = cell_4_7_out;
  // (4, 7) -> (4, 6) (out)
  assign cell_4_6_out = cell_4_7_out;
  // (5, 7) -> (6, 7) (out)
  assign cell_6_7_out = cell_5_7_out;
  // (5, 7) -> (4, 7) (out)
  assign cell_4_7_out = cell_5_7_out;
  // (5, 7) -> (5, 8) (out)
  assign cell_5_8_out = cell_5_7_out;
  // (5, 7) -> (5, 6) (out)
  assign cell_5_6_out = cell_5_7_out;
  // (6, 7) -> (7, 7) (out)
  assign cell_7_7_out = cell_6_7_out;
  // (6, 7) -> (5, 7) (out)
  assign cell_5_7_out = cell_6_7_out;
  // (6, 7) -> (6, 8) (out)
  assign cell_6_8_out = cell_6_7_out;
  // (6, 7) -> (6, 6) (out)
  assign cell_6_6_out = cell_6_7_out;
  // (7, 7) -> (8, 7) (out)
  assign cell_8_7_out = cell_7_7_out;
  // (7, 7) -> (6, 7) (out)
  assign cell_6_7_out = cell_7_7_out;
  // (7, 7) -> (7, 8) (out)
  assign cell_7_8_out = cell_7_7_out;
  // (7, 7) -> (7, 6) (out)
  assign cell_7_6_out = cell_7_7_out;
  // (8, 7) -> (9, 7) (out)
  assign cell_9_7_out = cell_8_7_out;
  // (8, 7) -> (7, 7) (out)
  assign cell_7_7_out = cell_8_7_out;
  // (8, 7) -> (8, 8) (out)
  assign cell_8_8_out = cell_8_7_out;
  // (8, 7) -> (8, 6) (out)
  assign cell_8_6_out = cell_8_7_out;
  // (9, 7) -> (10, 7) (out)
  assign cell_10_7_out = cell_9_7_out;
  // (9, 7) -> (8, 7) (out)
  assign cell_8_7_out = cell_9_7_out;
  // (9, 7) -> (9, 8) (out)
  assign cell_9_8_out = cell_9_7_out;
  // (9, 7) -> (9, 6) (out)
  assign cell_9_6_out = cell_9_7_out;
  // (10, 7) -> (11, 7) (out)
  assign cell_11_7_out = cell_10_7_out;
  // (10, 7) -> (9, 7) (out)
  assign cell_9_7_out = cell_10_7_out;
  // (10, 7) -> (10, 8) (out)
  assign cell_10_8_out = cell_10_7_out;
  // (10, 7) -> (10, 6) (out)
  assign cell_10_6_out = cell_10_7_out;
  // (11, 7) -> (10, 7) (out)
  assign cell_10_7_out = cell_11_7_out;
  // (11, 7) -> (11, 8) (out)
  assign cell_11_8_out = cell_11_7_out;
  // (11, 7) -> (11, 6) (out)
  assign cell_11_6_out = cell_11_7_out;
  // (0, 8) -> (1, 8) (out)
  assign cell_1_8_out = cell_0_8_out;
  // (0, 8) -> (0, 9) (out)
  assign cell_0_9_out = cell_0_8_out;
  // (0, 8) -> (0, 7) (out)
  assign cell_0_7_out = cell_0_8_out;
  // (1, 8) -> (2, 8) (out)
  assign cell_2_8_out = cell_1_8_out;
  // (1, 8) -> (0, 8) (out)
  assign cell_0_8_out = cell_1_8_out;
  // (1, 8) -> (1, 9) (out)
  assign cell_1_9_out = cell_1_8_out;
  // (1, 8) -> (1, 7) (out)
  assign cell_1_7_out = cell_1_8_out;
  // (2, 8) -> (3, 8) (out)
  assign cell_3_8_out = cell_2_8_out;
  // (2, 8) -> (1, 8) (out)
  assign cell_1_8_out = cell_2_8_out;
  // (2, 8) -> (2, 9) (out)
  assign cell_2_9_out = cell_2_8_out;
  // (2, 8) -> (2, 7) (out)
  assign cell_2_7_out = cell_2_8_out;
  // (3, 8) -> (4, 8) (out)
  assign cell_4_8_out = cell_3_8_out;
  // (3, 8) -> (2, 8) (out)
  assign cell_2_8_out = cell_3_8_out;
  // (3, 8) -> (3, 9) (out)
  assign cell_3_9_out = cell_3_8_out;
  // (3, 8) -> (3, 7) (out)
  assign cell_3_7_out = cell_3_8_out;
  // (4, 8) -> (5, 8) (out)
  assign cell_5_8_out = cell_4_8_out;
  // (4, 8) -> (3, 8) (out)
  assign cell_3_8_out = cell_4_8_out;
  // (4, 8) -> (4, 9) (out)
  assign cell_4_9_out = cell_4_8_out;
  // (4, 8) -> (4, 7) (out)
  assign cell_4_7_out = cell_4_8_out;
  // (5, 8) -> (6, 8) (out)
  assign cell_6_8_out = cell_5_8_out;
  // (5, 8) -> (4, 8) (out)
  assign cell_4_8_out = cell_5_8_out;
  // (5, 8) -> (5, 9) (out)
  assign cell_5_9_out = cell_5_8_out;
  // (5, 8) -> (5, 7) (out)
  assign cell_5_7_out = cell_5_8_out;
  // (6, 8) -> (7, 8) (out)
  assign cell_7_8_out = cell_6_8_out;
  // (6, 8) -> (5, 8) (out)
  assign cell_5_8_out = cell_6_8_out;
  // (6, 8) -> (6, 9) (out)
  assign cell_6_9_out = cell_6_8_out;
  // (6, 8) -> (6, 7) (out)
  assign cell_6_7_out = cell_6_8_out;
  // (7, 8) -> (8, 8) (out)
  assign cell_8_8_out = cell_7_8_out;
  // (7, 8) -> (6, 8) (out)
  assign cell_6_8_out = cell_7_8_out;
  // (7, 8) -> (7, 9) (out)
  assign cell_7_9_out = cell_7_8_out;
  // (7, 8) -> (7, 7) (out)
  assign cell_7_7_out = cell_7_8_out;
  // (8, 8) -> (9, 8) (out)
  assign cell_9_8_out = cell_8_8_out;
  // (8, 8) -> (7, 8) (out)
  assign cell_7_8_out = cell_8_8_out;
  // (8, 8) -> (8, 9) (out)
  assign cell_8_9_out = cell_8_8_out;
  // (8, 8) -> (8, 7) (out)
  assign cell_8_7_out = cell_8_8_out;
  // (9, 8) -> (10, 8) (out)
  assign cell_10_8_out = cell_9_8_out;
  // (9, 8) -> (8, 8) (out)
  assign cell_8_8_out = cell_9_8_out;
  // (9, 8) -> (9, 9) (out)
  assign cell_9_9_out = cell_9_8_out;
  // (9, 8) -> (9, 7) (out)
  assign cell_9_7_out = cell_9_8_out;
  // (10, 8) -> (11, 8) (out)
  assign cell_11_8_out = cell_10_8_out;
  // (10, 8) -> (9, 8) (out)
  assign cell_9_8_out = cell_10_8_out;
  // (10, 8) -> (10, 9) (out)
  assign cell_10_9_out = cell_10_8_out;
  // (10, 8) -> (10, 7) (out)
  assign cell_10_7_out = cell_10_8_out;
  // (11, 8) -> (10, 8) (out)
  assign cell_10_8_out = cell_11_8_out;
  // (11, 8) -> (11, 9) (out)
  assign cell_11_9_out = cell_11_8_out;
  // (11, 8) -> (11, 7) (out)
  assign cell_11_7_out = cell_11_8_out;
  // (0, 9) -> (1, 9) (out)
  assign cell_1_9_out = cell_0_9_out;
  // (0, 9) -> (0, 10) (out)
  assign cell_0_10_out = cell_0_9_out;
  // (0, 9) -> (0, 8) (out)
  assign cell_0_8_out = cell_0_9_out;
  // (1, 9) -> (2, 9) (out)
  assign cell_2_9_out = cell_1_9_out;
  // (1, 9) -> (0, 9) (out)
  assign cell_0_9_out = cell_1_9_out;
  // (1, 9) -> (1, 10) (out)
  assign cell_1_10_out = cell_1_9_out;
  // (1, 9) -> (1, 8) (out)
  assign cell_1_8_out = cell_1_9_out;
  // (2, 9) -> (3, 9) (out)
  assign cell_3_9_out = cell_2_9_out;
  // (2, 9) -> (1, 9) (out)
  assign cell_1_9_out = cell_2_9_out;
  // (2, 9) -> (2, 10) (out)
  assign cell_2_10_out = cell_2_9_out;
  // (2, 9) -> (2, 8) (out)
  assign cell_2_8_out = cell_2_9_out;
  // (3, 9) -> (4, 9) (out)
  assign cell_4_9_out = cell_3_9_out;
  // (3, 9) -> (2, 9) (out)
  assign cell_2_9_out = cell_3_9_out;
  // (3, 9) -> (3, 10) (out)
  assign cell_3_10_out = cell_3_9_out;
  // (3, 9) -> (3, 8) (out)
  assign cell_3_8_out = cell_3_9_out;
  // (4, 9) -> (5, 9) (out)
  assign cell_5_9_out = cell_4_9_out;
  // (4, 9) -> (3, 9) (out)
  assign cell_3_9_out = cell_4_9_out;
  // (4, 9) -> (4, 10) (out)
  assign cell_4_10_out = cell_4_9_out;
  // (4, 9) -> (4, 8) (out)
  assign cell_4_8_out = cell_4_9_out;
  // (5, 9) -> (6, 9) (out)
  assign cell_6_9_out = cell_5_9_out;
  // (5, 9) -> (4, 9) (out)
  assign cell_4_9_out = cell_5_9_out;
  // (5, 9) -> (5, 10) (out)
  assign cell_5_10_out = cell_5_9_out;
  // (5, 9) -> (5, 8) (out)
  assign cell_5_8_out = cell_5_9_out;
  // (6, 9) -> (7, 9) (out)
  assign cell_7_9_out = cell_6_9_out;
  // (6, 9) -> (5, 9) (out)
  assign cell_5_9_out = cell_6_9_out;
  // (6, 9) -> (6, 10) (out)
  assign cell_6_10_out = cell_6_9_out;
  // (6, 9) -> (6, 8) (out)
  assign cell_6_8_out = cell_6_9_out;
  // (7, 9) -> (8, 9) (out)
  assign cell_8_9_out = cell_7_9_out;
  // (7, 9) -> (6, 9) (out)
  assign cell_6_9_out = cell_7_9_out;
  // (7, 9) -> (7, 10) (out)
  assign cell_7_10_out = cell_7_9_out;
  // (7, 9) -> (7, 8) (out)
  assign cell_7_8_out = cell_7_9_out;
  // (8, 9) -> (9, 9) (out)
  assign cell_9_9_out = cell_8_9_out;
  // (8, 9) -> (7, 9) (out)
  assign cell_7_9_out = cell_8_9_out;
  // (8, 9) -> (8, 10) (out)
  assign cell_8_10_out = cell_8_9_out;
  // (8, 9) -> (8, 8) (out)
  assign cell_8_8_out = cell_8_9_out;
  // (9, 9) -> (10, 9) (out)
  assign cell_10_9_out = cell_9_9_out;
  // (9, 9) -> (8, 9) (out)
  assign cell_8_9_out = cell_9_9_out;
  // (9, 9) -> (9, 10) (out)
  assign cell_9_10_out = cell_9_9_out;
  // (9, 9) -> (9, 8) (out)
  assign cell_9_8_out = cell_9_9_out;
  // (10, 9) -> (11, 9) (out)
  assign cell_11_9_out = cell_10_9_out;
  // (10, 9) -> (9, 9) (out)
  assign cell_9_9_out = cell_10_9_out;
  // (10, 9) -> (10, 10) (out)
  assign cell_10_10_out = cell_10_9_out;
  // (10, 9) -> (10, 8) (out)
  assign cell_10_8_out = cell_10_9_out;
  // (11, 9) -> (10, 9) (out)
  assign cell_10_9_out = cell_11_9_out;
  // (11, 9) -> (11, 10) (out)
  assign cell_11_10_out = cell_11_9_out;
  // (11, 9) -> (11, 8) (out)
  assign cell_11_8_out = cell_11_9_out;
  // (0, 10) -> (1, 10) (out)
  assign cell_1_10_out = cell_0_10_out;
  // (0, 10) -> (0, 11) (out)
  assign cell_0_11_out = cell_0_10_out;
  // (0, 10) -> (0, 9) (out)
  assign cell_0_9_out = cell_0_10_out;
  // (1, 10) -> (2, 10) (out)
  assign cell_2_10_out = cell_1_10_out;
  // (1, 10) -> (0, 10) (out)
  assign cell_0_10_out = cell_1_10_out;
  // (1, 10) -> (1, 11) (out)
  assign cell_1_11_out = cell_1_10_out;
  // (1, 10) -> (1, 9) (out)
  assign cell_1_9_out = cell_1_10_out;
  // (2, 10) -> (3, 10) (out)
  assign cell_3_10_out = cell_2_10_out;
  // (2, 10) -> (1, 10) (out)
  assign cell_1_10_out = cell_2_10_out;
  // (2, 10) -> (2, 11) (out)
  assign cell_2_11_out = cell_2_10_out;
  // (2, 10) -> (2, 9) (out)
  assign cell_2_9_out = cell_2_10_out;
  // (3, 10) -> (4, 10) (out)
  assign cell_4_10_out = cell_3_10_out;
  // (3, 10) -> (2, 10) (out)
  assign cell_2_10_out = cell_3_10_out;
  // (3, 10) -> (3, 11) (out)
  assign cell_3_11_out = cell_3_10_out;
  // (3, 10) -> (3, 9) (out)
  assign cell_3_9_out = cell_3_10_out;
  // (4, 10) -> (5, 10) (out)
  assign cell_5_10_out = cell_4_10_out;
  // (4, 10) -> (3, 10) (out)
  assign cell_3_10_out = cell_4_10_out;
  // (4, 10) -> (4, 11) (out)
  assign cell_4_11_out = cell_4_10_out;
  // (4, 10) -> (4, 9) (out)
  assign cell_4_9_out = cell_4_10_out;
  // (5, 10) -> (6, 10) (out)
  assign cell_6_10_out = cell_5_10_out;
  // (5, 10) -> (4, 10) (out)
  assign cell_4_10_out = cell_5_10_out;
  // (5, 10) -> (5, 11) (out)
  assign cell_5_11_out = cell_5_10_out;
  // (5, 10) -> (5, 9) (out)
  assign cell_5_9_out = cell_5_10_out;
  // (6, 10) -> (7, 10) (out)
  assign cell_7_10_out = cell_6_10_out;
  // (6, 10) -> (5, 10) (out)
  assign cell_5_10_out = cell_6_10_out;
  // (6, 10) -> (6, 11) (out)
  assign cell_6_11_out = cell_6_10_out;
  // (6, 10) -> (6, 9) (out)
  assign cell_6_9_out = cell_6_10_out;
  // (7, 10) -> (8, 10) (out)
  assign cell_8_10_out = cell_7_10_out;
  // (7, 10) -> (6, 10) (out)
  assign cell_6_10_out = cell_7_10_out;
  // (7, 10) -> (7, 11) (out)
  assign cell_7_11_out = cell_7_10_out;
  // (7, 10) -> (7, 9) (out)
  assign cell_7_9_out = cell_7_10_out;
  // (8, 10) -> (9, 10) (out)
  assign cell_9_10_out = cell_8_10_out;
  // (8, 10) -> (7, 10) (out)
  assign cell_7_10_out = cell_8_10_out;
  // (8, 10) -> (8, 11) (out)
  assign cell_8_11_out = cell_8_10_out;
  // (8, 10) -> (8, 9) (out)
  assign cell_8_9_out = cell_8_10_out;
  // (9, 10) -> (10, 10) (out)
  assign cell_10_10_out = cell_9_10_out;
  // (9, 10) -> (8, 10) (out)
  assign cell_8_10_out = cell_9_10_out;
  // (9, 10) -> (9, 11) (out)
  assign cell_9_11_out = cell_9_10_out;
  // (9, 10) -> (9, 9) (out)
  assign cell_9_9_out = cell_9_10_out;
  // (10, 10) -> (11, 10) (out)
  assign cell_11_10_out = cell_10_10_out;
  // (10, 10) -> (9, 10) (out)
  assign cell_9_10_out = cell_10_10_out;
  // (10, 10) -> (10, 11) (out)
  assign cell_10_11_out = cell_10_10_out;
  // (10, 10) -> (10, 9) (out)
  assign cell_10_9_out = cell_10_10_out;
  // (11, 10) -> (10, 10) (out)
  assign cell_10_10_out = cell_11_10_out;
  // (11, 10) -> (11, 11) (out)
  assign cell_11_11_out = cell_11_10_out;
  // (11, 10) -> (11, 9) (out)
  assign cell_11_9_out = cell_11_10_out;
  // (0, 11) -> (1, 11) (out)
  assign cell_1_11_out = cell_0_11_out;
  // (0, 11) -> (0, 10) (out)
  assign cell_0_10_out = cell_0_11_out;
  // (1, 11) -> (2, 11) (out)
  assign cell_2_11_out = cell_1_11_out;
  // (1, 11) -> (0, 11) (out)
  assign cell_0_11_out = cell_1_11_out;
  // (1, 11) -> (1, 10) (out)
  assign cell_1_10_out = cell_1_11_out;
  // (2, 11) -> (3, 11) (out)
  assign cell_3_11_out = cell_2_11_out;
  // (2, 11) -> (1, 11) (out)
  assign cell_1_11_out = cell_2_11_out;
  // (2, 11) -> (2, 10) (out)
  assign cell_2_10_out = cell_2_11_out;
  // (3, 11) -> (4, 11) (out)
  assign cell_4_11_out = cell_3_11_out;
  // (3, 11) -> (2, 11) (out)
  assign cell_2_11_out = cell_3_11_out;
  // (3, 11) -> (3, 10) (out)
  assign cell_3_10_out = cell_3_11_out;
  // (4, 11) -> (5, 11) (out)
  assign cell_5_11_out = cell_4_11_out;
  // (4, 11) -> (3, 11) (out)
  assign cell_3_11_out = cell_4_11_out;
  // (4, 11) -> (4, 10) (out)
  assign cell_4_10_out = cell_4_11_out;
  // (5, 11) -> (6, 11) (out)
  assign cell_6_11_out = cell_5_11_out;
  // (5, 11) -> (4, 11) (out)
  assign cell_4_11_out = cell_5_11_out;
  // (5, 11) -> (5, 10) (out)
  assign cell_5_10_out = cell_5_11_out;
  // (6, 11) -> (7, 11) (out)
  assign cell_7_11_out = cell_6_11_out;
  // (6, 11) -> (5, 11) (out)
  assign cell_5_11_out = cell_6_11_out;
  // (6, 11) -> (6, 10) (out)
  assign cell_6_10_out = cell_6_11_out;
  // (7, 11) -> (8, 11) (out)
  assign cell_8_11_out = cell_7_11_out;
  // (7, 11) -> (6, 11) (out)
  assign cell_6_11_out = cell_7_11_out;
  // (7, 11) -> (7, 10) (out)
  assign cell_7_10_out = cell_7_11_out;
  // (8, 11) -> (9, 11) (out)
  assign cell_9_11_out = cell_8_11_out;
  // (8, 11) -> (7, 11) (out)
  assign cell_7_11_out = cell_8_11_out;
  // (8, 11) -> (8, 10) (out)
  assign cell_8_10_out = cell_8_11_out;
  // (9, 11) -> (10, 11) (out)
  assign cell_10_11_out = cell_9_11_out;
  // (9, 11) -> (8, 11) (out)
  assign cell_8_11_out = cell_9_11_out;
  // (9, 11) -> (9, 10) (out)
  assign cell_9_10_out = cell_9_11_out;
  // (10, 11) -> (11, 11) (out)
  assign cell_11_11_out = cell_10_11_out;
  // (10, 11) -> (9, 11) (out)
  assign cell_9_11_out = cell_10_11_out;
  // (10, 11) -> (10, 10) (out)
  assign cell_10_10_out = cell_10_11_out;
  // (11, 11) -> (10, 11) (out)
  assign cell_10_11_out = cell_11_11_out;
  // (11, 11) -> (11, 10) (out)
  assign cell_11_10_out = cell_11_11_out;
endmodule